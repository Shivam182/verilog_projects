module FIR_filter();




endmodule
